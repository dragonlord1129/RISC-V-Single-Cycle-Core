module instruction_memory (
    input rst,
    input [31:0] A,

    output [31:0] RD
);
    reg [31:0] memory [1023:0];
    
endmodule